library verilog;
use verilog.vl_types.all;
entity Modulo_IN_mas_Modulo_Estado_vlg_vec_tst is
end Modulo_IN_mas_Modulo_Estado_vlg_vec_tst;
