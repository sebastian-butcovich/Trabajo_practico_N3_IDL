library verilog;
use verilog.vl_types.all;
entity Maquina_de_estado_TP2_vlg_sample_tst is
    port(
        pin_name1       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Maquina_de_estado_TP2_vlg_sample_tst;
