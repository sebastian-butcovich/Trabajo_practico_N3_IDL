library verilog;
use verilog.vl_types.all;
entity Maquina_de_estados_V2_TP3_vlg_sample_tst is
    port(
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Maquina_de_estados_V2_TP3_vlg_sample_tst;
