library verilog;
use verilog.vl_types.all;
entity Modulo_IN_mas_Modulo_Estado_vlg_check_tst is
    port(
        aux             : in     vl_logic;
        Memoria_01      : in     vl_logic;
        Memoria_02      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Modulo_IN_mas_Modulo_Estado_vlg_check_tst;
