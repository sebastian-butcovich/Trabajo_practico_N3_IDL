library verilog;
use verilog.vl_types.all;
entity Maquina_de_estado_TP2_vlg_vec_tst is
end Maquina_de_estado_TP2_vlg_vec_tst;
