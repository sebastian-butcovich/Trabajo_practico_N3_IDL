library verilog;
use verilog.vl_types.all;
entity Trabajo_practico_03_Entrada_in_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        P0              : in     vl_logic;
        P1              : in     vl_logic;
        P2              : in     vl_logic;
        P3              : in     vl_logic;
        P4              : in     vl_logic;
        P5              : in     vl_logic;
        P6              : in     vl_logic;
        P7              : in     vl_logic;
        P8              : in     vl_logic;
        P9              : in     vl_logic;
        P10             : in     vl_logic;
        P11             : in     vl_logic;
        P12             : in     vl_logic;
        P13             : in     vl_logic;
        P14             : in     vl_logic;
        P15             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Trabajo_practico_03_Entrada_in_vlg_sample_tst;
