library verilog;
use verilog.vl_types.all;
entity Maquina_de_estados_V2_TP3_vlg_vec_tst is
end Maquina_de_estados_V2_TP3_vlg_vec_tst;
