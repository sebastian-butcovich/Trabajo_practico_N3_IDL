library verilog;
use verilog.vl_types.all;
entity Trabajo_practico_03_Entrada_in is
    port(
        S8              : out    vl_logic;
        CLK             : in     vl_logic;
        P8              : in     vl_logic;
        S9              : out    vl_logic;
        P9              : in     vl_logic;
        S10             : out    vl_logic;
        P10             : in     vl_logic;
        S11             : out    vl_logic;
        P11             : in     vl_logic;
        S12             : out    vl_logic;
        P12             : in     vl_logic;
        S13             : out    vl_logic;
        P13             : in     vl_logic;
        S14             : out    vl_logic;
        P14             : in     vl_logic;
        S15             : out    vl_logic;
        P15             : in     vl_logic;
        S7              : out    vl_logic;
        P7              : in     vl_logic;
        S6              : out    vl_logic;
        P6              : in     vl_logic;
        S5              : out    vl_logic;
        P5              : in     vl_logic;
        S4              : out    vl_logic;
        P4              : in     vl_logic;
        S3              : out    vl_logic;
        P3              : in     vl_logic;
        S2              : out    vl_logic;
        P2              : in     vl_logic;
        S1              : out    vl_logic;
        P1              : in     vl_logic;
        S0              : out    vl_logic;
        P0              : in     vl_logic
    );
end Trabajo_practico_03_Entrada_in;
