library verilog;
use verilog.vl_types.all;
entity Paralele_serie_16bits_vlg_check_tst is
    port(
        Salida          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Paralele_serie_16bits_vlg_check_tst;
