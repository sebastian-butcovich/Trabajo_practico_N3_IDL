library verilog;
use verilog.vl_types.all;
entity Paralele_serie_16bits_vlg_vec_tst is
end Paralele_serie_16bits_vlg_vec_tst;
